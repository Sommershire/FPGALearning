module tb_counter();



endmodule